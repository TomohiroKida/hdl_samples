module a();
endmodule
